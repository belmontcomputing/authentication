module hello;
endmodule
