module abc;
endmodule
