module v1;
endmodule
