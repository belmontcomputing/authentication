module v2;
endmodule
