module my_repo;
endmodule
