module my_repo_2;
endmodule
